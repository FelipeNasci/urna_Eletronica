library verilog;
use verilog.vl_types.all;
entity urna_vlg_vec_tst is
end urna_vlg_vec_tst;
